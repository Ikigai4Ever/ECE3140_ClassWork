--      Name: Ty Ahrens
--      Date: 10/31/2023
--      Purpose: VGA controller for DE10-Lite board

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity hw7p1 is 
    port(SW : IN std_logic_vector(2 downto 0);
         color_out : std_logic_vector(2 downto 0));
end hw7p1;




architecture Behavioral of hw7p1 is

end Behavioral;
