--Name: Ty Ahrens 
--Date: 3/30/2025
--Purpose: 

library IEEE;
use IEEE.std_logic_1164.all;

entity hw6 is 
    port();
end hw6;

architecture behavior of hw6 is 



end behavior;